// Code your testbench here
// or browse Examples
`include "apb_top.sv"
